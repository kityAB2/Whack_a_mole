module vga_display(
    input             vga_clk,                  //VGA驱动时钟
    input             sys_rst_n,                //复位信号
    input      [1:0]  page,                     //指示当前需要显示的页面
	input             mode,                     //指示当前显示的模式
	input      [3:0]  state,                     //指示当前需要显示的页面
	input      [3:0]  m,						//随机数
    input      [ 10:0] pixel_xpos,               //像素点横坐标
    input      [ 10:0] pixel_ypos,               //像素点纵坐标    
    output reg [23:0] pixel_data                //像素点数据,
    );    

//parameter define    
parameter  H_DISP = 11'd800;                    //分辨率——行
parameter  V_DISP = 11'd600;                    //分辨率——列
parameter INIT_ST = 4'd0;//游戏过程中状态机显示格子
parameter PIC1_ST = 4'd1;//游戏过程中状态机显示地鼠
parameter PIC2_ST = 4'd2;//游戏过程中状态机显示地鼠
parameter LINE_WIDTH = 11'd5;//网格线宽

localparam TITLE_POS_X  = 11'd48;                    //标题字符起始位置X
localparam TITLE_POS_Y  = 11'd80;                    //标题字符起始位置Y
localparam TITLE_WIDTH  = 11'd704;                     //字符区域宽度
localparam TITLE_HEIGHT = 11'd64;                     //字符区域高度

localparam MODE1_POS_X  = 11'd272;                    //标题字符起始位置X
localparam MODE1_POS_Y  = 11'd250;                    //标题字符起始位置Y
localparam MODE1_WIDTH  = 11'd256;                     //字符区域宽度
localparam MODE1_HEIGHT = 11'd64;                     //字符区域高度

localparam MODE2_POS_X  = 11'd272;                    //标题字符起始位置X
localparam MODE2_POS_Y  = 11'd350;                    //标题字符起始位置Y
localparam MODE2_WIDTH  = 11'd256;                     //字符区域宽度
localparam MODE2_HEIGHT = 11'd64;                     //字符区域高度
//游戏结束显示
localparam OVER_POS_X  = 11'd208;                    //标题字符起始位置X
localparam OVER_POS_Y  = 11'd270;                    //标题字符起始位置Y
localparam OVER_WIDTH  = 11'd384;                     //字符区域宽度
localparam OVER_HEIGHT = 11'd64;                     //字符区域高度
//游戏图片显示
//localparam POS_X  = 10'd270;                //图片区域起始点横坐标
//localparam POS_Y  = 10'd190;                //图片区域起始点纵坐标
localparam PIC1_WIDTH  = 11'd130;                //图片区域宽度
localparam PIC1_HEIGHT = 11'd130;                //图片区域高度
localparam PIC2_WIDTH  = 11'd130;                //图片区域宽度
localparam PIC2_HEIGHT = 11'd130;                //图片区域高度
localparam TOTAL  = 15'd16900;              //图案区域总像素数
reg [10:0] POS_X;                //图片区域起始点横坐标
reg [10:0] POS_Y;                //图片区域起始点纵坐标
//reg define rom1
wire        rom1_rd_en;                      //读ROM1使能信号
reg  [14:0] rom1_addr;                       //读ROM1地址
reg         rom1_valid;                      //读ROM1数据有效信号  
wire [23:0] rom1_data;                       //ROM1输出数据

//reg define rom2
wire        rom2_rd_en;                      //读ROM2使能信号
reg  [14:0] rom2_addr;                       //读ROM2地址
reg         rom2_valid;                      //读ROM2数据有效信号  
wire [23:0] rom2_data;                       //ROM2输出数据

localparam RED    = 24'b11111111_00000000_00000000;     //字符颜色
localparam BLUE   = 24'b00000000_00000000_11111111;     //字符区域背景色
localparam BLACK  = 24'b00000000_00000000_00000000;     //屏幕背景色
localparam WHITE  = 24'b11111111_11111111_11111111;     //白色

//reg define
reg  [703:0] title_char[63:0];                         //字符数组  
wire [ 10:0] title_x_cnt;
wire [ 10:0] title_y_cnt;
reg  [255:0] mode1_char[63:0];                         //字符数组  
wire [ 10:0] mode1_x_cnt;
wire [ 10:0] mode1_y_cnt;
reg  [255:0] mode2_char[63:0];                         //字符数组  
wire [ 10:0] mode2_x_cnt;
wire [ 10:0] mode2_y_cnt;
reg  [383:0] over_char[63:0];                         //字符数组  
wire [ 10:0] over_x_cnt;
wire [ 10:0] over_y_cnt;
//*****************************************************
//**                    main code
//*****************************************************
assign title_x_cnt = pixel_xpos - TITLE_POS_X;              //标题像素点相对于字符区域起始点水平坐标
assign title_y_cnt = pixel_ypos - TITLE_POS_Y;              //标题像素点相对于字符区域起始点竖直坐标
assign mode1_x_cnt = pixel_xpos - MODE1_POS_X;              //标题像素点相对于字符区域起始点水平坐标
assign mode1_y_cnt = pixel_ypos - MODE1_POS_Y;              //标题像素点相对于字符区域起始点竖直坐标
assign mode2_x_cnt = pixel_xpos - MODE2_POS_X;              //标题像素点相对于字符区域起始点水平坐标
assign mode2_y_cnt = pixel_ypos - MODE2_POS_Y;              //标题像素点相对于字符区域起始点竖直坐标
assign over_x_cnt = pixel_xpos - OVER_POS_X;              //标题像素点相对于字符区域起始点水平坐标
assign over_y_cnt = pixel_ypos - OVER_POS_Y;              //标题像素点相对于字符区域起始点竖直坐标
//给字符数组赋值，显示汉字“游戏难度选择”，汉字大小为64*64
always @(posedge vga_clk) begin
    title_char[0]  <= 704'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    title_char[1]  <= 704'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    title_char[2]  <= 704'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000600000000000000000000000000000000000000000000000000000000;
    title_char[3]  <= 704'h00000000000000000000800000000000000000000100000000000080000000000000000000100000000000004000000000000000004000000000000380000000000000000400000000010000000000000000000000000000;
    title_char[4]  <= 704'h00000000000000000000E000000000000000000001C00000000001C00000800000000000001C00000000000078000000000000001830000000000001E000000000000000070000000001C000000000000000000000000000;
    title_char[5]  <= 704'h00000001FFFFFE000000F80000000000000C000001F00000000007E00001C00000C00300001F0000000000007E000000000000003E38000000000001F00000000000000007C000000001F80000000800007FFFFF00000000;
    title_char[6]  <= 704'h00000001FFFFFC000000F00000000000000F000001E0000000001FF0FFFFE00000700180003E0000000000007E000000000000003F1C000000000000F80000000040000007C000000001F00000001C00003FFFFF00000000;
    title_char[7]  <= 704'h00000001FFFFF8000000E00000000000000F800001C000000018FF807FFFF000007C01E0003C0000000000007C000000000000003E1F0000000000007800030000300000070000000001E03FFFFFFE00001FFFFF00000000;
    title_char[8]  <= 704'h00000001FFFFF0000000E00000000080000F000001C00000001FF0002001E000003E00F000380000000000007C1C0000000000003C0F000000200000780007800038000C070000000001E01FFFFFFF00000FFFFF00000000;
    title_char[9]  <= 704'h00000001FFFFF0000000E000000001C0000F000001C00000001E00000001C000001F007800780000000000003C0F800000000000780F00000030000030000FC0001C000E070000000001E00080003E000007FFFF00000000;
    title_char[10] <= 704'h00000001FFFFE0000000E000000003E0000F000001C00000001E00000001C000001F007C00700000000000003C07E0000000000078070000003FFFFFFFFFFFE0001E001F870000000001E000400078000003FFFF00000000;
    title_char[11] <= 704'h00000001FFFFC0000000E00FFFFFFFF0000F000801C00000001E00000001C000000F003C00700080000000003C03F0000000010078070000003FFFFFFFFFFFF0000F001E070000000001E0006000F8000003FFFF00000000;
    title_char[12] <= 704'h00000001FFFF80000000E007FFFFFFF8000F000E01C00000001E00000001C000000F003800E00180000000003C01F800000001C070070000003C000000000000000F001E070000000001E0006000F0000001FFFF00000000;
    title_char[13] <= 704'h00000001FFFF80000000E000001E0000000F000F81C00000001E00600001C0000006003800E003C0000001803C00FC0007FFFFE0F0060300003C004000000000000F801C070000000001E0003001E0000000FFFF00000000;
    title_char[14] <= 704'h00000001FFFF00000000E060001E0000000F000F01C00000001E00F00001C0000000000001FFFFE0000003C03C007C0003FFFFF0E0000780003C0030001800000007801C070060000001E0003003C0000000FFFF00000000;
    title_char[15] <= 704'h00000001FFFE00000000E0F0001E0000000F000E01C00000001FFFF07FFFC0000000000081FFFFF00FFFFFE03C003800010003E0FFFFFFC0003C003C001E0000000780380700F0000001E0601807800000007FFF00000000;
	title_char[16] <= 704'h00000001FFFE00001FFFFFF8001E0000000F000E01C00800001FFFF83FFFC00000002001C180000007FFFFE03C003800000003C1FFFFFFE0003C003C001F00000007003FFFFFF8000001E0F00C0F800000007FFF00000000;
    title_char[17] <= 704'h00000001FFFC00000FFFFFFC001E0000000F000E01C01C00001E00001801C00000007FFFE3000000020007C01C00100000000381E01E0000003C0038001C00000002003FFFFFFC001FFFFFF80E1F000000003FFF00000000;
    title_char[18] <= 704'h00000001FFFC00000400E000001E0000000F000E01C03E00001E00000001C00010005FFFF3000000000007801C00018000000781E01E0000003C0038001C020000000070070000000FFFFFFC073E000000001FFF00000000;
    title_char[19] <= 704'h00000001FFF800000000E000001E0000000F000E01C0FF00001E00000001C0001C004DC006000000000007801E0001C000000783E01E0000003C0038001C070000000060070000000601E00007FC000000001FFF00000000;
    title_char[20] <= 704'h00000001FFF800000000E000001E0000000F000E01C3DE00001E00000001C0000F00C1C00C000100000007801E0003E000000783E01E0000003C0038001C0F80000000E0070000000001E00003F8000000001FFF00000000;
    title_char[21] <= 704'h00000001FFF000000000E000001E0000000F000E01CF1C00001E00000001C000078081C008000380000007801E000FF003000703E01E0000003FFFFFFFFFFFC0000000C0070000000001E00001F0000000000FFF00000000;
    title_char[22] <= 704'h00000001FFF000000000E000001E0000000F0C0E01F81C00001FFFFFFFFFC00007C081C013FFFFC000000F001E1FFFC001800F07E01E0000003DFFFFFFFFFFE0000000C0070000000001E00003F8000000000FFF00000000;
    title_char[23] <= 704'h00000001FFF000000000E000001E0000000F1E0E01C01C00001FFFFFFFFFC00003E181C011FFFFE000000F003FFF000000800F07E01E0000003C0038001C000000000180070000000001E00007FE0000000007FF00000000;
    title_char[24] <= 704'h00000001FFE000000000E000001E00001FFFFF0E0FC01C00001E00000001E00003E181C000C007C002000FFFFE00000000C00E0FE01E0000003C0038001C000000020300070000000001E0001F1FC000000007FF00000000;
    title_char[25] <= 704'h00000001FFE000000000E000001E00000FFFFF8E79C01C00001E00000001000001E101C000000F0003000E7C0E00000000600E0FE01E0000003C0038001C000000070200070006000001E0103C0FF800000007FF00000000;
    title_char[26] <= 704'h00000001FFE000000000E018001E0000040F000FE1C01C00001000080000000001E301C060001C0001801E200F00000000301E1DE01E0600003C0038001C00001FFF800007000F000001E060F903FFF8000007FF00000000;
    title_char[27] <= 704'h00000001FFE000000000E0F0001E0000000F001F01C01C000000000E0008000000C301FFF000380000E01E000F00080000181C19E01E0F00003C0038001C00000FFF9FFFFFFFFF800001E1C1E1C0FFF0000003FF00000000;
    title_char[28] <= 704'h00000001FFE000000000E3C0001E0000000F007E01C01C000010000F800E0000008301FFF800600000701E000F001C00001C1C39FFFFFF80003C0038001C0000040F0FFFFFFFFFC00001E70781F03FC0000003FF00000000;
    title_char[29] <= 704'h00000001FFC000000000EF00001E0000000F03CE01C01C00001C000F800F0000000201C0F002400000381C000F001E00000E3C31FFFFFFC000380038001C0000000F0400E07800000001FE1E01F80F80000003FF00000000;
    title_char[30] <= 704'h00000001FFC000000000FC00001E0000000F1E0E01C01C00001F700F200F0000000601C0E0038000001C3C000F003F0000073861E01E00000038003FFFFC0000000F0000E07800000001F87801E00100000003FF00000000;
    title_char[31] <= 704'h00000001FFC000000003F000001E0000000F1C0E01C01C00001E3C0F380E0000000601C0E003E000000E3C0007003E0000073841E01E00000038003FFFFC0000000F0000E07800000003F1C001E00000000003FF00000000;
	title_char[32] <= 704'h00000001FFC00000001FE000001E0000000F000E01C01C00001E1F0F1E0E0000000603C0E003C0000007380007807C000003F8C1E01E000000380038001C0000000F0001E0780000000FE30001E00000000003FF00000000;
	title_char[33] <= 704'h00000001FFC0000000FFE000001E0000000F000E01C01C00001E0F8F0F8E0000000C03C0E003C0000007F8000780F8000001F181E01E00000038003000180000000F0001E0780000007FE00001E00C00000003FF00000000;
    title_char[34] <= 704'h00000001FFC0000007FCE000001E0000000F000E01C01C00001E078F07CE0000000C0380E003C0000003F8000780F0000000F001E01E00000038004000010000000F0001E078000001FDE00001E01E00000003FF00000000;
    title_char[35] <= 704'h00000001FFC000000FF0E000001E0000000F000E01C01C00001E038F03CE0000000C0380E003C0C00001F0000381F0000000F001E01E00000078000000038000000F0001C07800000FF1E03FFFFFFF00000007FF00000000;
    title_char[36] <= 704'h00000001FFE0000007C0E000001E0000000F000E01C01C00001E038F01CE0000001C0380E003C1E00000F0000383E0000001F001E01E000000781FFFFFFFC000000F0001C07800000FE1E01FFFFFFF80000007FF00000000;
    title_char[37] <= 704'h00000001FFE000000380E000001E0000000F000E01C01C00001E018F01CF000000180380EFFFFFE00001F80003C7C0000001F801E01E020000780FFFFFFFE000000F0003C07800000F81E00801E00000000007FF00000000;
    title_char[38] <= 704'h00000001FFE000000200E000001E0000000F000E01C01C00001E000F008F000000380380E7FFFFF00001FC0003C780000003FC01E01E0700007000200007C000000F0003807801800701E00001E00000000007FF00000000;
    title_char[39] <= 704'h00000001FFE000000000E000001E0000000F000E01C01C00001E000F2007000000380700E203C0000003FE0001CF800000039E01E01E0F8000700010000F8000000F0003807801800201E00001E00000000007FF00000000;
    title_char[40] <= 704'h00000001FFF000000000E000001E0000000F000E01DFFC00001E700F3C07000000780700E003C00000039F0001FF000000079E01FFFFFFC000700018001F0000000F0007807801800001E00001E0000000000FFF00000000;
    title_char[41] <= 704'h00000001FFF000000000E000001E0000000F000E01C3FC00001E3C0F1F0700001FF00701C003C00000039F0001FE000000070F01FFFFFFE00070000C003E0000000F0007007801800001E00001E0000000000FFF00000000;
    title_char[42] <= 704'h00000001FFF000000000E000001E0000000F000E01C0F800001E1E0F0F87000007F00701C003C00000070F8000FC0020000E0F01E01E00000070000E003C0000000F000F007801800001E00001E0008000000FFF00000000;
    title_char[43] <= 704'h00000001FFF800000000E000001E0000000F000E01C07840001E1F0F0787000001F00E01C003C000000F07C000F80020001C0781E01E000000E0000700780000000F000E007801800001E00001E001C000001FFF00000000;
    title_char[44] <= 704'h00000001FFF800000000E000001E0000000F00CE01C02040001E0F0F03C7800000F00E01C003C000000E07C001F00020001C0781E01E000000E0000300F80000000F001C007801800001E00001E003E000001FFF00000000;
    title_char[45] <= 704'h00000001FFFC00000000E000001E0000000F078E01C00040001E070F0383804000F00E01C003C000001C03E003F8002000380381E01E000000E00001C1F00000000F0038007001800001E3FFFFFFFFF000003FFF00000000;
    title_char[46] <= 704'h00000001FFFC00000000E000001E0000000F3E0E01C00040001E070F0183804000F01C01C003C000001C03E007FC0020007003C1E01E000000E00001E3E00000000F0070007803800001E1FFFFFFFFF800003FFF00000000;
    title_char[47] <= 704'h00000001FFFE00000000E000001E0000000FF80E01800040001E020F018380C000F01C01C003C000003801E00FBE0060006003C1E01E000000C00000F7C00000000F00E0007803E00001E0C001E0000000007FFF00000000;
	title_char[48] <= 704'h00000001FFFE00000000E000001E0000000FC00E02000040001E000F0003C0C000F03801C003C000003001E01F1E006000C003C1E01E000001C000007F800000001F01C0003FFFE00001E00001E0000000007FFF00000000;
    title_char[49] <= 704'h00000001FFFF00000000E000001E0000007F000E00000060001E010F0101C08001F03803C003C000007000C03C0F006001C00181E01E0000018000003F000000007F8380003FFFC00001E00001E000000000FFFF00000000;
    title_char[50] <= 704'h00000001FFFF80000000E000001E000003FC000E000000E0001E070F0601E18001E070038003C00000E000C0780F806003800181E01E0000018000003E00000001F1CE00001FFF800001E00001E000000001FFFF00000000;
    title_char[51] <= 704'h00000001FFFF80000000E000001E00003FF0000E000000E0001E1C0F3C00F18001E070038003C00000C00000F007C0E007000001E01E000003800000FF80000003E0E800000000000001E00001E000000001FFFF00000000;
    title_char[52] <= 704'h00000001FFFFC0000000E000001E00001FC0000E000000F0001E780FF800F18001E0E0038003C00001800003C003F0E006000001E01E00C003000001FFE000000FC03800000000000001E00001E000000003FFFF00000000;
    title_char[53] <= 704'h00000001FFFFE0000201E000001E00000F80000E000000F8001FE00FE0007B8001E0C0078003C000038000078001F8E008000001E01E01E003000007E3FC00001F801C00000000000001E00001E000000007FFFF00000000;
    title_char[54] <= 704'h00000001FFFFE00003FBE0007E3C00000E00000F000001F8001FC00FC0003F8001E183FF8003C0000700000E0000FEE010000001FFFFFFF00600001F80FF80003F000F800000000003C3E00001E000000007FFFF00000000;
    title_char[55] <= 704'h00000001FFFFF00000FFE0001FFC00000400000FFFFFFFF0003F800F80003F8000E380FF01FFC0000600003800007FE000000001FFFFFFF80600007E007FFE000E0007FE000003FC01FFE00001E00000000FFFFF00000000;
    title_char[56] <= 704'h00000001FFFFF800003FE00007FC000000000007FFFFFFF0001F000700001F800063007E007FC0000C00007000003FE000000001E00000000C0003F0001FFFF0060001FFFFFFFFE0003FC00001E00000001FFFFF00000000;
    title_char[57] <= 704'h00000001FFFFFC00000FC00001F8000000000003FFFFFFC0000E000200000FC00006003E001F8000180001C000001FE000000001E000000008000FC00003FFC00000007FFFFFFFC0001FC00001E00000003FFFFF00000000;
    title_char[58] <= 704'h00000001FFFFFE000007C00000F80000000000000000000000040002000003C0000C0038000F800030000700000007F000000001E000000018007E0000007F8000000007FFFFFF80000F800001E00000007FFFFF00000000;
    title_char[59] <= 704'h00000000000000000003800000E00000000000000000000000000000000000C0001800000007000000000400000001F000000001E00000001007E00000000F000000000007FFFF000007000001E000000000000000000000;
    title_char[60] <= 704'h0000000000000000000200000000000000000000000000000000000000000000001000000000000000000000000000380000000100000000201C000000000000000000000000000000040000018000000000000000000000;
    title_char[61] <= 704'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    title_char[62] <= 704'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    title_char[63] <= 704'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	mode1_char[0]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    mode1_char[1]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    mode1_char[2]  <= 256'h0000000000000000000000000000000000000000004000000000000000000000;
    mode1_char[3]  <= 256'h0000000000000000000000000200000000003000006000000000000000000000;
    mode1_char[4]  <= 256'h0000000000000000000380000300000000001C00007800000000000000000000;
    mode1_char[5]  <= 256'h00000001FFFFFE000003C0000780000000000E0000FC0000007FFFFF00000000;
    mode1_char[6]  <= 256'h00000001FFFFFC000007E00007E000000000078000F80000003FFFFF00000000;
    mode1_char[7]  <= 256'h00000001FFFFF8000007C0000F800000000007C001F00000001FFFFF00000000;
    mode1_char[8]  <= 256'h00000001FFFFF000000F80080F000300000003E001E00000000FFFFF00000000;
    mode1_char[9]  <= 256'h00000001FFFFF000000F001C1E000780000003E001C000000007FFFF00000000;
    mode1_char[10] <= 256'h00000001FFFFE000001FFFFE1FFFFFC0000001E0038000000003FFFF00000000;
    mode1_char[11] <= 256'h00000001FFFFC000001FFFFFBFFFFFE0000001E0030000000003FFFF00000000;
    mode1_char[12] <= 256'h00000001FFFF80000038300078300000000000E0060000000001FFFF00000000;
    mode1_char[13] <= 256'h00000001FFFF800000701C00701C0000000800C00C0000000000FFFF00000000;
    mode1_char[14] <= 256'h00000001FFFF000000600E00E00E0000000C00000C00C0000000FFFF00000000;
    mode1_char[15] <= 256'h00000001FFFE000000C00F01C00F0000000FFFFFFFFFF00000007FFF00000000;
	mode1_char[16] <= 256'h00000001FFFE000001C00F01800F0000000FFFFFFFFFF00000007FFF00000000;
    mode1_char[17] <= 256'h00000001FFFC00000380070300070000000F00078001E00000003FFF00000000;
    mode1_char[18] <= 256'h00000001FFFC00000303070600060000000F00078001E00000001FFF00000000;
    mode1_char[19] <= 256'h00000001FFF800000403800400000000000F00078001E00000001FFF00000000;
    mode1_char[20] <= 256'h00000001FFF800000801E00000000C00000F00078001E00000001FFF00000000;
    mode1_char[21] <= 256'h00000001FFF000000000F07FFFFFFE00000F00078001E00000000FFF00000000;
    mode1_char[22] <= 256'h00000001FFF000000000783FFFFFFF00000F00078001E00000000FFF00000000;
    mode1_char[23] <= 256'h00000001FFF0000000407C1000001E00000F00078001E000000007FF00000000;
    mode1_char[24] <= 256'h00000001FFE0000000303C0000001C00000FFFFFFFFFE000000007FF00000000;
    mode1_char[25] <= 256'h00000001FFE00000003C3C0000001C00000FFFFFFFFFE000000007FF00000000;
    mode1_char[26] <= 256'h00000001FFE00000003C380000001C00000F00078001E000000007FF00000000;
    mode1_char[27] <= 256'h00000001FFE000000038100000001C00000F00078001E000000003FF00000000;
    mode1_char[28] <= 256'h00000001FFE000000038000002001C00000F00078001E000000003FF00000000;
    mode1_char[29] <= 256'h00000001FFC000000038018003001C00000F00078001E000000003FF00000000;
    mode1_char[30] <= 256'h00000001FFC00000003801FFFF801C00000F00078001E000000003FF00000000;
    mode1_char[31] <= 256'h00000001FFC00000003801FFFFC01C00000F00078001E000000003FF00000000;
	mode1_char[32] <= 256'h00000001FFC00000003801E007801C00000F00078001E000000003FF00000000;
	mode1_char[33] <= 256'h00000001FFC00000003801E007001C00000F00078001E000000003FF00000000;
    mode1_char[34] <= 256'h00000001FFC00000003801E007001C00000FFFFFFFFFE000000003FF00000000;
    mode1_char[35] <= 256'h00000001FFC00000003801E007001C00000FFFFFFFFFE000000007FF00000000;
    mode1_char[36] <= 256'h00000001FFE00000003801E007001C00000F00078001E000000007FF00000000;
    mode1_char[37] <= 256'h00000001FFE00000003801E007001C00000F00078001C000000007FF00000000;
    mode1_char[38] <= 256'h00000001FFE00000003801E007001C00000F000780010000000007FF00000000;
    mode1_char[39] <= 256'h00000001FFE00000003801FFFF001C00000E000780000000000007FF00000000;
    mode1_char[40] <= 256'h00000001FFF00000003801FFFF001C00000000078000000000000FFF00000000;
    mode1_char[41] <= 256'h00000001FFF00000003801E007001C00000000078000018000000FFF00000000;
    mode1_char[42] <= 256'h00000001FFF00000003801E007001C0000000007800003C000000FFF00000000;
    mode1_char[43] <= 256'h00000001FFF80000003801E007001C0000000007800007E000001FFF00000000;
    mode1_char[44] <= 256'h00000001FFF80000003801E007001C001FFFFFFFFFFFFFF000001FFF00000000;
    mode1_char[45] <= 256'h00000001FFFC0000003801E007001C000FFFFFFFFFFFFFF800003FFF00000000;
    mode1_char[46] <= 256'h00000001FFFC0000003801E007001C00000000078000000000003FFF00000000;
    mode1_char[47] <= 256'h00000001FFFE0000003801E007001C00000000078000000000007FFF00000000;
	mode1_char[48] <= 256'h00000001FFFE0000003801FFFF001C00000000078000000000007FFF00000000;
    mode1_char[49] <= 256'h00000001FFFF0000003801FFFF001C0000000007800000000000FFFF00000000;
    mode1_char[50] <= 256'h00000001FFFF8000003801E007001C0000000007800000000001FFFF00000000;
    mode1_char[51] <= 256'h00000001FFFF8000003801E006001C0000000007800000000001FFFF00000000;
    mode1_char[52] <= 256'h00000001FFFFC000003801E000001C0000000007800000000003FFFF00000000;
    mode1_char[53] <= 256'h00000001FFFFE0000038010000001C0000000007800000000007FFFF00000000;
    mode1_char[54] <= 256'h00000001FFFFE0000038000000001C0000000007800000000007FFFF00000000;
    mode1_char[55] <= 256'h00000001FFFFF00000380000007C3C000000000780000000000FFFFF00000000;
    mode1_char[56] <= 256'h00000001FFFFF80000380000001FFC000000000780000000001FFFFF00000000;
    mode1_char[57] <= 256'h00000001FFFFFC00003800000003FC000000000780000000003FFFFF00000000;
    mode1_char[58] <= 256'h00000001FFFFFE00003800000001FC000000000780000000007FFFFF00000000;
    mode1_char[59] <= 256'h0000000000000000003800000000780000000007800000000000000000000000;
    mode1_char[60] <= 256'h0000000000000000003800000000600000000004000000000000000000000000;
    mode1_char[61] <= 256'h0000000000000000002000000000000000000000000000000000000000000000;
    mode1_char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
    mode1_char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	mode2_char[0]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;		
	mode2_char[1]  <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	mode2_char[2]  <= 256'h0000000000000000000000000000000000000000040000000000000000000000;
	mode2_char[3]  <= 256'h0000000000000000000000010008000000000000070000000000000000000000;
	mode2_char[4]  <= 256'h000000000000000000000001C00E0000000000000F8000000000000000000000;
	mode2_char[5]  <= 256'h00000001FFFFFE0000400001F00F8000040008000F800000007FFFFF00000000;
	mode2_char[6]  <= 256'h00000001FFFFFC0000300001F00F800006001C000F000000003FFFFF00000000;
	mode2_char[7]  <= 256'h00000001FFFFF800003C0001E00F000007FFFE001F800000001FFFFF00000000;
	mode2_char[8]  <= 256'h00000001FFFFF000001E0001C00F000007FFFF001E800000000FFFFF00000000;
	mode2_char[9]  <= 256'h00000001FFFFF000000F0001C00F000007803E003CC000000007FFFF00000000;
	mode2_char[10] <= 256'h00000001FFFFE000000F8001C00F000007803C003C6000000003FFFF00000000;
	mode2_char[11] <= 256'h00000001FFFFC00000078001C00F000007807800786000000003FFFF00000000;
	mode2_char[12] <= 256'h00000001FFFF80000007C001C00F000007807800703000000001FFFF00000000;
	mode2_char[13] <= 256'h00000001FFFF800000078001C00F020007807000F03800000000FFFF00000000;
	mode2_char[14] <= 256'h00000001FFFF000000038001C00F060007807000E01C00000000FFFF00000000;
	mode2_char[15] <= 256'h00000001FFFE000000030001C00F0F000780E001C01C000000007FFF00000000;
	mode2_char[16] <= 256'h00000001FFFE000000000FFFFFFFFF800780E003C00E000000007FFF00000000;
	mode2_char[17] <= 256'h00000001FFFC0000000007FFFFFFFFC00780C0078007000000003FFF00000000;
	mode2_char[18] <= 256'h00000001FFFC000000000301C00F00000781C0070007C00000001FFF00000000;
	mode2_char[19] <= 256'h00000001FFF8000000000001C00F00000781800E0003E00000001FFF00000000;
	mode2_char[20] <= 256'h00000001FFF8000000000001C00F00000781801C0001F80000001FFF00000000;
	mode2_char[21] <= 256'h00000001FFF0000000000001C00F0000078300380000FE0000000FFF00000000;
	mode2_char[22] <= 256'h00000001FFF0000000000001C00F00000783007000007F8000000FFF00000000;
	mode2_char[23] <= 256'h00000001FFF0000000020001C00F0000078200E000001FF0000007FF00000000;
	mode2_char[24] <= 256'h00000001FFE0000000070001C00F0000078601C000080FF8000007FF00000000;
	mode2_char[25] <= 256'h00000001FFE000003FFF8001C00F000007830301000E07E0000007FF00000000;
	mode2_char[26] <= 256'h00000001FFE000001FFFC001C00F000007818601C00F01C0000007FF00000000;
	mode2_char[27] <= 256'h00000001FFE00000080F0001C00F00000780C801F00F8000000003FF00000000;
	mode2_char[28] <= 256'h00000001FFE00000000F0001C00F000007804001C00F0000000003FF00000000;
	mode2_char[29] <= 256'h00000001FFC00000000F0001C00F000007806001C00F0000000003FF00000000;
	mode2_char[30] <= 256'h00000001FFC00000000F0001C00F018007803001C00F0000000003FF00000000;
	mode2_char[31] <= 256'h00000001FFC00000000F0001C00F03C007803801C00F0000000003FF00000000;
	mode2_char[32] <= 256'h00000001FFC00000000F1FFFFFFFFFE007803801C00F0000000003FF00000000;
	mode2_char[33] <= 256'h00000001FFC00000000F0FFFFFFFFFF007801C01C00F0000000003FF00000000;
	mode2_char[34] <= 256'h00000001FFC00000000F0401C00F000007801C01C00F0000000003FF00000000;
	mode2_char[35] <= 256'h00000001FFC00000000F0001C00F000007801C01C00F0000000007FF00000000;
	mode2_char[36] <= 256'h00000001FFE00000000F0001C00F000007801E01C00F0000000007FF00000000;
	mode2_char[37] <= 256'h00000001FFE00000000F0001C00F000007801E01C00F0000000007FF00000000;
	mode2_char[38] <= 256'h00000001FFE00000000F0003800F000007801E01C00F0000000007FF00000000;
	mode2_char[39] <= 256'h00000001FFE00000000F0003800F000007801E01C00F0000000007FF00000000;
	mode2_char[40] <= 256'h00000001FFF00000000F0003800F000007803C03C00F000000000FFF00000000;
	mode2_char[41] <= 256'h00000001FFF00000000F0007000F000007F87C03C00F000000000FFF00000000;
	mode2_char[42] <= 256'h00000001FFF00000000F0007000F000007FFFC03C00F000000000FFF00000000;
	mode2_char[43] <= 256'h00000001FFF80000000F000E000F0000079FF803800F000000001FFF00000000;
	mode2_char[44] <= 256'h00000001FFF80000000F000E000F00000787F003800F000000001FFF00000000;
	mode2_char[45] <= 256'h00000001FFFC0000000F001C000F00000783E003800F000000003FFF00000000;
	mode2_char[46] <= 256'h00000001FFFC0000000F0038000F000007838003800F000000003FFF00000000;
	mode2_char[47] <= 256'h00000001FFFE0000000F0070000F000007800007800F000000007FFF00000000;
	mode2_char[48] <= 256'h00000001FFFE0000000F00E0000F000007800007000F000000007FFF00000000;
	mode2_char[49] <= 256'h00000001FFFF0000001F81C0000F000007800007000F00000000FFFF00000000;
	mode2_char[50] <= 256'h00000001FFFF80000039C300000F00000780000E000F00000001FFFF00000000;
	mode2_char[51] <= 256'h00000001FFFF80000070E400000F00000780000E000F00000001FFFF00000000;
	mode2_char[52] <= 256'h00000001FFFFC00001E03800000E00000780001C000F00000003FFFF00000000;
	mode2_char[53] <= 256'h00000001FFFFE00003C01E000008000007800018000F00000007FFFF00000000;
	mode2_char[54] <= 256'h00000001FFFFE00007800F800000000007800038000F00000007FFFF00000000;
	mode2_char[55] <= 256'h00000001FFFFF0000F8007FC0000007C07800070000F0000000FFFFF00000000;
	mode2_char[56] <= 256'h00000001FFFFF8001F0001FFFFFFFFF0078000C0000F0000001FFFFF00000000;
	mode2_char[57] <= 256'h00000001FFFFFC000E00007FFFFFFFC007800180000F0000003FFFFF00000000;
	mode2_char[58] <= 256'h00000001FFFFFE000600001FFFFFFF8007800700000E0000007FFFFF00000000;
	mode2_char[59] <= 256'h0000000000000000000000003FFFFF0007000C00000800000000000000000000;
	mode2_char[60] <= 256'h0000000000000000000000000000000004001000000000000000000000000000;
	mode2_char[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	mode2_char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	mode2_char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	over_char[0]  <= 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;	
	over_char[1]  <= 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	over_char[2]  <= 384'h000000000000000000000000000000000000000000000000000000000080000000000002000000000000000000000000;
	over_char[3]  <= 384'h0000000000000000000000000010000000000000400000000001000000E0000000000003800000000000000000000000;
	over_char[4]  <= 384'h000000000000000000000000001C000000000000780000000001C00000F8000000000003E00000000000000000000000;
	over_char[5]  <= 384'h00000000FFFFFE0000C00300001F0000000000007E0000000001F00000FC000000000003E0000000007FFFFF00000000;
	over_char[6]  <= 384'h00000000FFFFFC0000700180003E0000000000007E0000000003F00000F0000000000003C0000000003FFFFF00000000;
	over_char[7]  <= 384'h00000000FFFFF800007C01E0003C0000000000007C0000000003C00000F0000000000003C0000000001FFFFF00000000;
	over_char[8]  <= 384'h00000000FFFFF000003E00F000380000000000007C1C00000003C00000F0000000000003C0000100000FFFFF00000000;	
	over_char[9]  <= 384'h00000000FFFFE000001F007800780000000000003C0F80000007800000F0000000000003C00003800007FFFF00000000;
	over_char[10] <= 384'h00000000FFFFC000001F007C00700000000000003C07E0000007800000F0000000000003C00007C00003FFFF00000000;
	over_char[11] <= 384'h00000000FFFFC000000F003C00700080000000003C03F0000007000000F000000FFFFFFFFFFFFFE00003FFFF00000000;
	over_char[12] <= 384'h00000000FFFF8000000F003800E00180000000003C01F800000E000000F0000007FFFFFFFFFFFFF00001FFFF00000000;
	over_char[13] <= 384'h00000000FFFF00000006003800E003C0000001803C00FC00000E000000F0018002000003C00000000000FFFF00000000;
	over_char[14] <= 384'h00000000FFFF00000000000001FFFFE0000003C03C007C00001C000000F003C000000003C00000000000FFFF00000000;
	over_char[15] <= 384'h00000000FFFE00000000000081FFFFF00FFFFFE03C003800001C003FFFFFFFE000000003C000000000007FFF00000000;
	over_char[16] <= 384'h00000000FFFE000000002001C180000007FFFFE03C0038000018001FFFFFFFF000000003C000000000007FFF00000000;	
	over_char[17] <= 384'h00000000FFFC000000007FFFE3000000020007C01C0010000038038800F0000000000003C000000000003FFF00000000;
	over_char[18] <= 384'h00000000FFF8000010005FFFF3000000000007801C000180003003C000F0000000000003C000C00000001FFF00000000;
	over_char[19] <= 384'h00000000FFF800001C004DC006000000000007801E0001C0006007E000F00000000C0003C000E00000001FFF00000000;
	over_char[20] <= 384'h00000000FFF800000F00C1C00C000100000007801E0003E00060078000F00000000FFFFFFFFFF80000001FFF00000000;
	over_char[21] <= 384'h00000000FFF00000078081C008000380000007801E000FF000C00F0000F00000000FFFFFFFFFF80000000FFF00000000;
	over_char[22] <= 384'h00000000FFF0000007C081C013FFFFC000000F001E1FFFC001C01F0000F00000000F0003C001E00000000FFF00000000;
	over_char[23] <= 384'h00000000FFE0000003E181C011FFFFE000000F003FFF000001801E0000F00000000F0003C001E000000007FF00000000;
	over_char[24] <= 384'h00000000FFE0000003E181C000C007C002000FFFFE00000003003C0000F00000000F0003C001E000000007FF00000000;	
	over_char[25] <= 384'h00000000FFE0000001E101C000000F0003000E7C0E0000000FFFF80000F00400000F0003C001E000000007FF00000000;
	over_char[26] <= 384'h00000000FFE0000001E301C060001C0001801E200F00000007FFF00000F00C00000F0003C001E000000007FF00000000;
	over_char[27] <= 384'h00000000FFC0000000C301FFF000380000E01E000F00080007F0F00000F01E00000F0003C001E000000003FF00000000;
	over_char[28] <= 384'h00000000FFC00000008301FFF800600000701E000F001C000380E00FFFFFFF00000F0003C001E000000003FF00000000;
	over_char[29] <= 384'h00000000FFC00000000201C0F002400000381C000F001E000201C007FFFFFF80000F0003C001E000000003FF00000000;
	over_char[30] <= 384'h00000000FFC00000000601C0E0038000001C3C000F003F000003800300000000000F0003C001E000000003FF00000000;
	over_char[31] <= 384'h00000000FFC00000000601C0E003E000000E3C0007003E000003000000000000000F0003C001E000000003FF00000000;
	over_char[32] <= 384'h00000000FFC00000000603C0E003C0000007380007807C000007000000000000000F0003C001E000000003FF00000000;	
	over_char[33] <= 384'h00000000FFC00000000C03C0E003C0000007F8000780F800000E000000000000000F0003C001E000000003FF00000000;
	over_char[34] <= 384'h00000000FFC00000000C0380E003C0000003F8000780F000001C000000000000000FFFFFFFFFE000000003FF00000000;
	over_char[35] <= 384'h00000000FFC00000000C0380E003C0C00001F0000381F0000038000200000400000FFFFFFFFFE000000007FF00000000;
	over_char[36] <= 384'h00000000FFC00000001C0380E003C1E00000F0000383E0000030000300000E00000F003FD001E000000007FF00000000;
	over_char[37] <= 384'h00000000FFE0000000180380EFFFFFE00001F80003C7C00000600FE3FFFFFF00000F007FD801E000000007FF00000000;
	over_char[38] <= 384'h00000000FFE0000000380380E7FFFFF00001FC0003C7800001C3FE03FFFFFF80000F007BC801C000000007FF00000000;
	over_char[39] <= 384'h00000000FFE0000000380700E203C0000003FE0001CF800003FFF003C0001F00000F00FBCC010000000007FF00000000;
	over_char[40] <= 384'h00000000FFE0000000780700E003C00000039F0001FF000003FF0003C0001E00000C01F3C600000000000FFF00000000;	
	over_char[41] <= 384'h00000000FFF000001FF00701C003C00000039F0001FE000003F80003C0001E00000001E3C700000000000FFF00000000;
	over_char[42] <= 384'h00000000FFF0000007F00701C003C00000070F8000FC002001E00003C0001E00000003E3C300000000000FFF00000000;
	over_char[43] <= 384'h00000000FFF0000001F00E01C003C000000F07C000F8002000800003C0001E00000007C3C380000000001FFF00000000;
	over_char[44] <= 384'h00000000FFF8000000F00E01C003C000000E07C001F0002000000003C0001E0000000F83C1C0000000001FFF00000000;
	over_char[45] <= 384'h00000000FFF8000000F00E01C003C000001C03E003F8002000000003C0001E0000000F03C0E0000000003FFF00000000;
	over_char[46] <= 384'h00000000FFFC000000F01C01C003C000001C03E007FC002000000013C0001E0000001E03C070000000003FFF00000000;
	over_char[47] <= 384'h00000000FFFC000000F01C01C003C000003801E00FBE0060000000F3C0001E0000003C03C07C000000007FFF00000000;
	over_char[48] <= 384'h00000000FFFE000000F03801C003C000003001E01F1E006000000783C0001E0000007803C03E000000007FFF00000000;	
	over_char[49] <= 384'h00000000FFFF000001F03803C003C000007000C03C0F006000007E03C0001E000000F003C01F80000000FFFF00000000;
	over_char[50] <= 384'h00000000FFFF000001E070038003C00000E000C0780F80600003F803C0001E000001E003C00FC0000001FFFF00000000;
	over_char[51] <= 384'h00000000FFFF800001E070038003C00000C00000F007C0E0007FC003C0001E000003C003C007F0000001FFFF00000000;
	over_char[52] <= 384'h00000000FFFFC00001E0E0038003C00001800003C003F0E00FFF0003C0001E00000F8003C003FE000003FFFF00000000;
	over_char[53] <= 384'h00000000FFFFC00001E0C0078003C000038000078001F8E00FFC0003FFFFFE00001E0003C001FFC00007FFFF00000000;
	over_char[54] <= 384'h00000000FFFFE00001E183FF8003C0000700000E0000FEE007F00003FFFFFE00003C0003C0007FF00007FFFF00000000;
	over_char[55] <= 384'h00000000FFFFF00000E380FF01FFC0000600003800007FE007C00003C0001E0000700003C0003FC0000FFFFF00000000;
	over_char[56] <= 384'h00000000FFFFF8000063007E007FC0000C00007000003FE003000003C0001E0001E00003C0000F00001FFFFF00000000;	
	over_char[57] <= 384'h00000000FFFFFC000006003E001F8000180001C000001FE002000003C0001E0003800003C0000600003FFFFF00000000;
	over_char[58] <= 384'h00000000FFFFFE00000C0038000F800030000700000007F000000003C0001E000E000003C0000000007FFFFF00000000;
	over_char[59] <= 384'h0000000000000000001800000007000000000400000001F0000000038000180018000003C00000000000000000000000;
	over_char[60] <= 384'h000000000000000000100000000000000000000000000038000000020000000000000003800000000000000000000000;
	over_char[61] <= 384'h000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000;
	over_char[62] <= 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	over_char[63] <= 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end
//地址POs_X
always @(*) begin
    case (m)  
		4'b0000 : POS_X = 11'd35;
		4'b0001 : POS_X	= 11'd35+11'd200;
		4'b0010 : POS_X	= 11'd35+11'd200+11'd200;
		4'b0011 : POS_X	= 11'd35+11'd200+11'd200+11'd200;
		4'b0100 : POS_X	= 11'd35;
		4'b0101 : POS_X	= 11'd35+11'd200;	
		4'b0110 : POS_X	= 11'd35+11'd200+11'd200;
		4'b0111 : POS_X	= 11'd35+11'd200+11'd200+11'd200;
		4'b1000 : POS_X	= 11'd35;
		4'b1001 : POS_X	= 11'd35+11'd200;
		4'b1010 : POS_X	= 11'd35+11'd200+11'd200;
		4'b1011 : POS_X	= 11'd35+11'd200+11'd200+11'd200;
		4'b1100 : POS_X	= 11'd35;
		4'b1101 : POS_X	= 11'd35+11'd200;
		4'b1110 : POS_X	= 11'd35+11'd200+11'd200;
		4'b1111 : POS_X	= 11'd35+11'd200+11'd200+11'd200;
		default:;
	endcase 
end
//地址POs_Y
always @(*) begin
    case (m)  
		4'b0000 : POS_Y = 11'd10;
		4'b0001 : POS_Y	= 11'd10;
		4'b0010 : POS_Y	= 11'd10;
		4'b0011 : POS_Y	= 11'd10;
		4'b0100 : POS_Y	= 11'd10+11'd150;
		4'b0101 : POS_Y	= 11'd10+11'd150;	
		4'b0110 : POS_Y	= 11'd10+11'd150;
		4'b0111 : POS_Y	= 11'd10+11'd150;
		4'b1000 : POS_Y	= 11'd10+11'd150+11'd150;
		4'b1001 : POS_Y	= 11'd10+11'd150+11'd150;
		4'b1010 : POS_Y	= 11'd10+11'd150+11'd150;
		4'b1011 : POS_Y	= 11'd10+11'd150+11'd150;
		4'b1100 : POS_Y	= 11'd10+11'd150+11'd150+11'd150;
		4'b1101 : POS_Y	= 11'd10+11'd150+11'd150+11'd150;
		4'b1110 : POS_Y	= 11'd10+11'd150+11'd150+11'd150;
		4'b1111 : POS_Y	= 11'd10+11'd150+11'd150+11'd150;
		default:;  	
	endcase 
end
//给不同的区域绘制不同的颜色
always @(posedge vga_clk or negedge sys_rst_n) begin         
    if (!sys_rst_n) 
        pixel_data <= WHITE;
    else begin
		if(page==2'd0) begin//第一个界面
			if((pixel_xpos >= TITLE_POS_X) && (pixel_xpos < TITLE_POS_X + TITLE_WIDTH)//绘制标题
			  && (pixel_ypos >= TITLE_POS_Y) && (pixel_ypos < TITLE_POS_Y + TITLE_HEIGHT)) begin
				if(title_char[title_y_cnt][TITLE_WIDTH - title_x_cnt])
					pixel_data <= RED;              //绘制字符为红色
				else
					pixel_data <= WHITE;             //绘制字符区域背景为蓝色      
			end
			else if((pixel_xpos >= MODE1_POS_X) && (pixel_xpos < MODE1_POS_X + MODE1_WIDTH)//绘制模式
			  && (pixel_ypos >= MODE1_POS_Y) && (pixel_ypos < MODE1_POS_Y + MODE1_HEIGHT)) begin
				if(mode1_char[mode1_y_cnt][MODE1_WIDTH - mode1_x_cnt])
					pixel_data <= RED;              //绘制字符为红色
				else begin
					if(mode==1'b0) begin
						pixel_data <= BLUE;             //绘制字符区域背景为蓝色    
					end
					else pixel_data <= WHITE;             //绘制字符区域背景为白色 
				end
			end
			else if((pixel_xpos >= MODE2_POS_X) && (pixel_xpos < MODE2_POS_X + MODE2_WIDTH)//绘制模式
			  && (pixel_ypos >= MODE2_POS_Y) && (pixel_ypos < MODE2_POS_Y + MODE2_HEIGHT)) begin
				if(mode2_char[mode2_y_cnt][MODE2_WIDTH - mode2_x_cnt])
					pixel_data <= RED;              //绘制字符为红色
				else begin
					if(mode==1'b0) begin
						pixel_data <= WHITE;             //绘制字符区域背景为白色    
					end
					else pixel_data <= BLUE;             //绘制字符区域背景为蓝色
				end
			end
			else pixel_data <= WHITE;                //绘制屏幕背景为白色
		end
		else if(page==2'd1) begin//游戏模式
			if(state==INIT_ST) begin//绘制网格
				if((pixel_xpos>=11'd200-LINE_WIDTH) && (pixel_xpos<=11'd200+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_xpos>=11'd400-LINE_WIDTH) && (pixel_xpos<=11'd400+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_xpos>=11'd600-LINE_WIDTH) && (pixel_xpos<=11'd600+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_ypos>=11'd150-LINE_WIDTH) && (pixel_ypos<=11'd150+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_ypos>=11'd300-LINE_WIDTH) && (pixel_ypos<=11'd300+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_ypos>=11'd450-LINE_WIDTH) && (pixel_ypos<=11'd450+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else pixel_data <= WHITE;                //绘制屏幕背景为白色
			end
			else if(state==PIC1_ST) begin
				if((pixel_xpos>=11'd200-LINE_WIDTH) && (pixel_xpos<=11'd200+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_xpos>=11'd400-LINE_WIDTH) && (pixel_xpos<=11'd400+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_xpos>=11'd600-LINE_WIDTH) && (pixel_xpos<=11'd600+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_ypos>=11'd150-LINE_WIDTH) && (pixel_ypos<=11'd150+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_ypos>=11'd300-LINE_WIDTH) && (pixel_ypos<=11'd300+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_ypos>=11'd450-LINE_WIDTH) && (pixel_ypos<=11'd450+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_xpos >= POS_X) && (pixel_xpos < POS_X + PIC1_WIDTH)//显示对应的图片
						&& (pixel_ypos >= POS_Y) && (pixel_ypos < POS_Y + PIC1_HEIGHT)) begin
					pixel_data <= rom1_data;
			    end
				else pixel_data <= WHITE;                //绘制屏幕背景为白色
			end
			else if(state==PIC2_ST) begin
				if((pixel_xpos>=11'd200-LINE_WIDTH) && (pixel_xpos<=11'd200+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_xpos>=11'd400-LINE_WIDTH) && (pixel_xpos<=11'd400+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_xpos>=11'd600-LINE_WIDTH) && (pixel_xpos<=11'd600+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_ypos>=11'd150-LINE_WIDTH) && (pixel_ypos<=11'd150+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_ypos>=11'd300-LINE_WIDTH) && (pixel_ypos<=11'd300+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_ypos>=11'd450-LINE_WIDTH) && (pixel_ypos<=11'd450+LINE_WIDTH)) begin
					pixel_data <= RED;
				end
				else if((pixel_xpos >= POS_X) && (pixel_xpos < POS_X + PIC2_WIDTH)//显示对应的图片
						&& (pixel_ypos >= POS_Y) && (pixel_ypos < POS_Y + PIC2_HEIGHT)) begin
					pixel_data <= rom2_data;
			    end
				else pixel_data <= WHITE;                //绘制屏幕背景为白色
			
			end
		
		end
		else if(page==2'd2) begin//游戏结束模式
			if((pixel_xpos >= OVER_POS_X) && (pixel_xpos < OVER_POS_X + OVER_WIDTH)//绘制标题
			  && (pixel_ypos >= OVER_POS_Y) && (pixel_ypos < OVER_POS_Y + OVER_HEIGHT)) begin
				if(over_char[over_y_cnt][OVER_WIDTH - over_x_cnt])
					pixel_data <= RED;              //绘制字符为红色
				else
					pixel_data <= WHITE;             //绘制字符区域背景为蓝色      
			end
			
		end
    end
end
//assign pixel_data = rom_valid ? rom_data : BLACK; 
//当前像素点坐标位于图案显示区域内时，读ROM使能信号拉高
assign rom1_rd_en = (pixel_xpos >= POS_X-1'b1) && (pixel_xpos < POS_X + PIC1_WIDTH-1'b1)
                    && (pixel_ypos >= POS_Y) && (pixel_ypos < POS_Y + PIC1_HEIGHT)
                     ? 1'b1 : 1'b0;
//从发出读使能到ROM输出有效数据存在一个时钟周期的延时
//always @(posedge vga_clk or negedge sys_rst_n) begin         
//    if (!sys_rst_n) 
//        rom_valid <= 1'b0;
//    else
//        rom_valid <= rom_rd_en;
//end
//控制读地址
always @(posedge vga_clk or negedge sys_rst_n) begin         
    if (!sys_rst_n) begin
        rom1_addr   <= 15'd0;
    end
	else if(pixel_xpos==11'd1&&pixel_ypos==11'd1) begin
		rom1_addr   <= 15'd0;
	end
    else if(rom1_rd_en) begin
        if(rom1_addr < TOTAL - 1'b1)
            rom1_addr <= rom1_addr + 1'b1;    //每次读ROM操作后，读地址加1
        else
            rom1_addr <= 1'b0;               //读到ROM末地址后，从首地址重新开始读操作
    end
    else
        rom1_addr <= rom1_addr;
end
//通过调用IP核来例化ROM1
pic1_rom	pic1_rom_inst(
	.clock   (vga_clk),
	.address (rom1_addr),
	.rden    (rom1_rd_en),
	.q       (rom1_data)
	);
	
	
//assign pixel_data = rom_valid ? rom_data : BLACK; 
//当前像素点坐标位于图案显示区域内时，读ROM使能信号拉高
assign rom2_rd_en = (pixel_xpos >= POS_X-1'b1) && (pixel_xpos < POS_X + PIC2_WIDTH-1'b1)
                    && (pixel_ypos >= POS_Y) && (pixel_ypos < POS_Y + PIC2_HEIGHT)
                     ? 1'b1 : 1'b0;
//从发出读使能到ROM输出有效数据存在一个时钟周期的延时
//always @(posedge vga_clk or negedge sys_rst_n) begin         
//    if (!sys_rst_n) 
//        rom_valid <= 1'b0;
//    else
//        rom_valid <= rom_rd_en;
//end
//控制读地址
always @(posedge vga_clk or negedge sys_rst_n) begin         
    if (!sys_rst_n) begin
        rom2_addr   <= 15'd0;
    end
	else if(pixel_xpos==11'd1&&pixel_ypos==11'd1) begin
		rom2_addr   <= 15'd0;
	end
    else if(rom2_rd_en) begin
        if(rom2_addr < TOTAL - 1'b1)
            rom2_addr <= rom2_addr + 1'b1;    //每次读ROM操作后，读地址加1
        else
            rom2_addr <= 1'b0;               //读到ROM末地址后，从首地址重新开始读操作
    end
	else
		rom2_addr <= rom2_addr;
end
     	
//通过调用IP核来例化ROM2
pic2_rom	pic2_rom_inst(
	.clock   (vga_clk),
	.address (rom2_addr),
	.rden    (rom2_rd_en),
	.q       (rom2_data)
	);
endmodule 