module seg7(
    input     [3:0]          d    ,          // 数据输入
    input                    rst_n   ,       // 使能信号  低电平使能
    output    reg [6:0]      seg_data        // 
    );   
always @ (*)//组合电路
begin
    if(!rst_n) begin	        //判断使能
		seg_data[6:0] = ~(7'b0000000);					//判断输入的BCD码
    end
    else begin
		case (d)  
            4'b0000 : seg_data[6:0] = ~(7'b0111111);	//数码管将会显示 "0"
            4'b0001 : seg_data[6:0] = ~(7'b0000110);	//数码管将会显示 "1"
            4'b0010 : seg_data[6:0] = ~(7'b1011011);	//数码管将会显示 "2"
            4'b0011 : seg_data[6:0] = ~(7'b1001111);	//数码管将会显示 "3"
            4'b0100 : seg_data[6:0] = ~(7'b1100110);	//数码管将会显示 "4"
            4'b0101 : seg_data[6:0] = ~(7'b1101101);	//数码管将会显示 "5"	
            4'b0110 : seg_data[6:0] = ~(7'b1111101);	//数码管将会显示 "0"
            4'b0111 : seg_data[6:0] = ~(7'b0000111);	//数码管将会显示 "7"
            4'b1000 : seg_data[6:0] = ~(7'b1111111);	//数码管将会显示 "8"
            4'b1001 : seg_data[6:0] = ~(7'b1101111);	//数码管将会显示 "9"
            4'b1010 : seg_data[6:0] = ~(7'b1110111);	//数码管将会显示 "A"
            4'b1011 : seg_data[6:0] = ~(7'b1111100);	//数码管将会显示 "b"
            4'b1100 : seg_data[6:0] = ~(7'b0111001);	//数码管将会显示 "c"
            4'b1101 : seg_data[6:0] = ~(7'b1011110);	//数码管将会显示 "d"
            4'b1110 : seg_data[6:0] = ~(7'b1111001);	//数码管将会显示 "E"
            4'b1111 : seg_data[6:0] = ~(7'b1110001);	//数码管将会显示 "F"
		default:  seg_data[6:0] = ~(7'b0000000);	
	endcase 	
    end
end
endmodule